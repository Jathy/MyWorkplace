`timescale 1ns/1ps
//**********************************************************************
// 	Project: 
//	File: xxx.v
// 	Description: 
//	Author: Noa
//  Timestamp: 
//----------------------------------------------------------------------
// Code Revision History:
// Ver:		| Author 	| Mod. Date		| Changes Made:
// v1.0.0	| Noa		| xx/xx/20xx	| Initial version
//**********************************************************************
//`include "./define/define.vh"
module tb;

//**********************************************************************
// --- Parameter
//**********************************************************************
// `include "./define/parameter.vh"

	localparam CLK_PERIOD = 50.0;			
	localparam NUM_DATA = 20; 

//**********************************************************************
// --- Test Input signal
//**********************************************************************	
	reg 		sym_clk;
	reg			rstn;
	reg	[9:0]	data_reg;
	reg [9:0]	mem_data [0:21] = {50, 75, 100, 150, 196, 238, 271, 292, 300, 292, 271, 238, 196, 150, 103,  61,  28,  28,  61, 103, 149, 195};
	
/*
x = 0:2*pi/20:2*pi
y = floor(150*(sin(x)+1))  
 150   196   238   271   292   300   292   271   238   196   150   103    61 
    28     7     0     7    28    61   103   149
*/
//**********************************************************************
// --- Test Output signal
//**********************************************************************
	wire [9:0] data_event_intr;
	
//**********************************************************************
// --- Internal Signal Declaration
//**********************************************************************	

	

//**********************************************************************
// --- Define Variable	
//**********************************************************************	
	integer i_data;
	
//**********************************************************************	
// --- Initial Block
//**********************************************************************

	GSR GSR(.GSRI(1'b1));

	adc_event_ctrl adc_event_ctrl_inst(
		.adc_wclk		(sym_clk),
		.adc_wclk_rstn	(rstn),
		.data_reg		( data_reg),
		.data_v1_reg	( 10'd50 ),
		.data_v2_reg	( 10'd100 ),
		.data_v3_reg	( 10'd225 ),
		.data_v4_reg	( 10'd275 ),
		.data_v5_reg	( 10'd275 ),
		.data_v6_reg	( 10'd275 ),
		.data_v7_reg	( 10'd200 ),
		.data_v8_reg	( 10'd50 ),
		.data_v9_reg	( 10'd50 ),
		.data_v10_reg	( 10'd100 ),
		.data_event_en	( 10'b11_1111_1111),
		.data_event_mask( 10'b00_0000_0000),
		.data_event_intr( data_event_intr)
);

//**********************************************************************	
// --- Clock Generate
//**********************************************************************
	initial begin
		sym_clk = 1'b1;
		#(1.5*CLK_PERIOD) 
		forever #(CLK_PERIOD/2.0) sym_clk = ~sym_clk;
	end

//**********************************************************************
// --- Reset 
//**********************************************************************
	initial begin
		rstn = 1'b1;
		#(1.5*CLK_PERIOD) rstn = 1'b0;
		#(CLK_PERIOD) rstn = 1'b1;
	end
//**********************************************************************
// --- Constant Setting
//**********************************************************************



//**********************************************************************
// --- Read file
//**********************************************************************

//**********************************************************************
// --- Input simulation
//**********************************************************************
	initial begin
		data_reg = 0;
		
		#(3*CLK_PERIOD);
		
		for (i_data=0; i_data < NUM_DATA; i_data = i_data+1) begin
			#(CLK_PERIOD*10);
			data_reg = mem_data[i_data];
		end
		
		#(CLK_PERIOD*10);
	end
	

	
//**********************************************************************
// --- Write file
//**********************************************************************	
	// always @(posedge sym_clk) begin
		// if(sel_valid) $fdisplay(fid_wr,"%d",fir_data_d);
	// end

	// initial begin
        // fid_wr = $fopen(FILE_RESULT, "w");
        // $fsdbDumpfile("fir_tb.fsdb");
        // $fsdbDumpvars;
	// end
//**********************************************************************
// --- 
//**********************************************************************	
	// initial begin
		
	// end
	
endmodule
